Library ieee;
USE ieee.std_logic_1164.all;


ENTITY O_1 IS
PORT ( SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END O_1;

ARCHITECTURE Behavior OF O_1 IS
BEGIN
LEDR <= SW;
END Behavior;