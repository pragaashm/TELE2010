LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;


ENTITY O_3 IS
	PORT( 
	SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
	LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END O_3;

ARCHITECTURE muxUVWX OF O_3 IS
	SIGNAL U,V,W,X,Y : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL M : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL S : STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN

	S <= SW(9 DOWNTO 8);
	U <= SW(7 DOWNTO 6);
	V <= SW(5 DOWNTO 4);
	W <= SW(3 DOWNTO 2);
	X <= SW(1 DOWNTO 0);
	M <= (((NOT S(1) AND NOT S(0) AND U(0)) OR (NOT S(1) AND S(0) AND V(0)) OR (S(1) AND NOT S(0) AND W(0)) OR (S(1) AND S(0) AND X(0))), ((NOT S(1) AND NOT S(0) AND U(1)) OR (NOT S(1) AND S(0) AND V(1)) OR (S(1) AND NOT S(0) AND W(1)) OR (S(1) AND S(0) AND X(1)))); 
	LEDR(1 DOWNTO 0) <= M;	
	LEDR(9 DOWNTO 8) <= S;
	
	
END muxUVWX;